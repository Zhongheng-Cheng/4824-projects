
// P1 TODO: create the testbench. Use ps4_test as a starting point
