
module ps4 (
    input        [3:0] req,
    input              en,
    output logic [3:0] gnt
);

    // P1 TODO: use assign statements and logic to create a priority selector
    // do not use any always blocks
    // ex:
    // assign x = y[1] & z & ~a;


endmodule
