
module ISR (
    input               reset,
    input        [63:0] value,
    input               clock,
    output logic [31:0] result,
    output logic        done
);

    // P2 TODO: Finish answering questions for the mult module,
    //          then implement the Integer Square Root algorithm as specified

    // P2 NOTE: reset mult_defs.svh to 8 stages when using this module.

endmodule
